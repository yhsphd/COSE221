// AND Gate
module and2(x, y, s);

input x, y;
output s;

// RTL M
assign s=x&y;

endmodule 